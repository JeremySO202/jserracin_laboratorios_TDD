
`ifndef CONNECT4_TYPES_SV
`define CONNECT4_TYPES_SV

package connect4_tipos;


typedef enum logic [4:0] {
	INICIO,          
	MENU,
	JUGADOR_INICIAL,
	TURNO_J1,   // Turno del jugador 1 (FPGA)
	VERIFICAR_J1,
	TIEMPO_J1,
	RANDOM_J1,
	GANADOR_J1,
	FIN_JUEGO_J1,
	TURNO_J2,   // Turno del jugador 2 (Arduino)
	VERIFICAR_J2,
	TIEMPO_J2,
	RANDOM_J2,
	GANADOR_J2,
	FIN_JUEGO_J2
} game_state;

endpackage

`endif // CONNECT4_TYPES_SV