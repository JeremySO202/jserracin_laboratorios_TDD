`include "connect4_tipos.sv"

module connect4_fsm(
	input clk, rst, inicio_juego, num_jugador,
	input t_J1, valido_J1, gano_J1, tiempo_terminado_J1, random_valido_J1,
	input t_J2, valido_J2, gano_J2, tiempo_terminado_J2, random_valido_J2,
	output logic jugador, 
	output logic enTurno1, enTurno2, 
	output logic enVerificar1, enVerificar2, 
	output logic enGanador, 
	output logic finJuego1, finJuego2 
	);
	

	import connect4_tipos::*;
	logic [4:0] state, next_state;

//actual state

always_ff @(posedge clk or posedge rst)
	if (rst) state = INICIO;
	else
		state = next_state;


always_comb
	case(state)
	INICIO: next_state = MENU;
	MENU: next_state = inicio_juego? JUGADOR_INICIAL : MENU;
	JUGADOR_INICIAL: next_state = num_jugador? TURNO_J2 : TURNO_J1;
	TURNO_J1: next_state = t_J1? VERIFICAR_J1 : TIEMPO_J1;
	TIEMPO_J1: next_state = tiempo_terminado_J1? RANDOM_J1 : TURNO_J1;
	RANDOM_J1: next_state = random_valido_J1? GANADOR_J1 : RANDOM_J1;
	VERIFICAR_J1: next_state = valido_J1? GANADOR_J1 : TURNO_J1;
	GANADOR_J1: next_state = gano_J1? FIN_JUEGO_J1 : TURNO_J2;
	FIN_JUEGO_J1: next_state = FIN_JUEGO_J1;
	TURNO_J2: next_state = t_J2? VERIFICAR_J2 : TIEMPO_J2;
	TIEMPO_J2: next_state = tiempo_terminado_J2? RANDOM_J2 : TURNO_J2;
	RANDOM_J2: next_state = random_valido_J2? GANADOR_J2 : RANDOM_J2;
	VERIFICAR_J2: next_state = valido_J2? GANADOR_J2 : TURNO_J2;
	GANADOR_J2: next_state = gano_J2? FIN_JUEGO_J2 : TURNO_J1;
	FIN_JUEGO_J2: next_state = FIN_JUEGO_J2;
	default: next_state = INICIO;
	endcase

	assign jugador = (state == TURNO_J2) || (state == TIEMPO_J2) || (state == RANDOM_J2) || (state == VERIFICAR_J2) || (state == GANADOR_J2) || (state == FIN_JUEGO_J2); // Habilitar el turno del jugador 2
	
	assign enTurno1 = (state == TURNO_J1); // Habilitar el turno del jugador 1
	assign enVerificar1 = (state == VERIFICAR_J1); // Habilitar la verificación del jugador 1
	
	assign enTurno2 = (state == TURNO_J2); // Habilitar el turno del jugador 2
	assign enVerificar2 = (state == VERIFICAR_J2); // Habilitar la verificación del jugador 2

	assign enGanador = (state == GANADOR_J1) || (state == GANADOR_J2); // Habilitar la verificación del ganador

	assign finJuego1 = (state == FIN_JUEGO_J1); // Habilitar la verificación del jugador 1
	assign finJuego2 = (state == FIN_JUEGO_J2); // Habilitar la verificación del jugador 2

	
endmodule